##
## LEF for PtnCells ;
## created by Innovus v18.10-p002_1 on Fri Apr  2 20:41:29 2021
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO aes128key
  CLASS BLOCK ;
  SIZE 236.930000 BY 234.920000 ;
  FOREIGN aes128key -118.465000 -117.460000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 19.820000 234.850000 19.890000 234.920000 ;
    END
  END reset
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 20.580000 234.850000 20.650000 234.920000 ;
    END
  END clock
  PIN empty
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 21.340000 234.850000 21.410000 234.920000 ;
    END
  END empty
  PIN load
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 22.100000 234.850000 22.170000 234.920000 ;
    END
  END load
  PIN key[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 119.380000 234.850000 119.450000 234.920000 ;
    END
  END key[127]
  PIN key[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 118.620000 234.850000 118.690000 234.920000 ;
    END
  END key[126]
  PIN key[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 117.860000 234.850000 117.930000 234.920000 ;
    END
  END key[125]
  PIN key[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 117.100000 234.850000 117.170000 234.920000 ;
    END
  END key[124]
  PIN key[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 116.340000 234.850000 116.410000 234.920000 ;
    END
  END key[123]
  PIN key[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 115.580000 234.850000 115.650000 234.920000 ;
    END
  END key[122]
  PIN key[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 114.820000 234.850000 114.890000 234.920000 ;
    END
  END key[121]
  PIN key[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 114.060000 234.850000 114.130000 234.920000 ;
    END
  END key[120]
  PIN key[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 113.300000 234.850000 113.370000 234.920000 ;
    END
  END key[119]
  PIN key[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 112.540000 234.850000 112.610000 234.920000 ;
    END
  END key[118]
  PIN key[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 111.780000 234.850000 111.850000 234.920000 ;
    END
  END key[117]
  PIN key[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 111.020000 234.850000 111.090000 234.920000 ;
    END
  END key[116]
  PIN key[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 110.260000 234.850000 110.330000 234.920000 ;
    END
  END key[115]
  PIN key[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 109.500000 234.850000 109.570000 234.920000 ;
    END
  END key[114]
  PIN key[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 108.740000 234.850000 108.810000 234.920000 ;
    END
  END key[113]
  PIN key[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 107.980000 234.850000 108.050000 234.920000 ;
    END
  END key[112]
  PIN key[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 107.220000 234.850000 107.290000 234.920000 ;
    END
  END key[111]
  PIN key[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 106.460000 234.850000 106.530000 234.920000 ;
    END
  END key[110]
  PIN key[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 105.700000 234.850000 105.770000 234.920000 ;
    END
  END key[109]
  PIN key[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 104.940000 234.850000 105.010000 234.920000 ;
    END
  END key[108]
  PIN key[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 104.180000 234.850000 104.250000 234.920000 ;
    END
  END key[107]
  PIN key[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 103.420000 234.850000 103.490000 234.920000 ;
    END
  END key[106]
  PIN key[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 102.660000 234.850000 102.730000 234.920000 ;
    END
  END key[105]
  PIN key[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 101.900000 234.850000 101.970000 234.920000 ;
    END
  END key[104]
  PIN key[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 101.140000 234.850000 101.210000 234.920000 ;
    END
  END key[103]
  PIN key[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 100.380000 234.850000 100.450000 234.920000 ;
    END
  END key[102]
  PIN key[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 99.620000 234.850000 99.690000 234.920000 ;
    END
  END key[101]
  PIN key[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 98.860000 234.850000 98.930000 234.920000 ;
    END
  END key[100]
  PIN key[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 98.100000 234.850000 98.170000 234.920000 ;
    END
  END key[99]
  PIN key[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 97.340000 234.850000 97.410000 234.920000 ;
    END
  END key[98]
  PIN key[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 96.580000 234.850000 96.650000 234.920000 ;
    END
  END key[97]
  PIN key[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 95.820000 234.850000 95.890000 234.920000 ;
    END
  END key[96]
  PIN key[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 95.060000 234.850000 95.130000 234.920000 ;
    END
  END key[95]
  PIN key[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 94.300000 234.850000 94.370000 234.920000 ;
    END
  END key[94]
  PIN key[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 93.540000 234.850000 93.610000 234.920000 ;
    END
  END key[93]
  PIN key[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 92.780000 234.850000 92.850000 234.920000 ;
    END
  END key[92]
  PIN key[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 92.020000 234.850000 92.090000 234.920000 ;
    END
  END key[91]
  PIN key[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 91.260000 234.850000 91.330000 234.920000 ;
    END
  END key[90]
  PIN key[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 90.500000 234.850000 90.570000 234.920000 ;
    END
  END key[89]
  PIN key[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 89.740000 234.850000 89.810000 234.920000 ;
    END
  END key[88]
  PIN key[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 88.980000 234.850000 89.050000 234.920000 ;
    END
  END key[87]
  PIN key[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 88.220000 234.850000 88.290000 234.920000 ;
    END
  END key[86]
  PIN key[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 87.460000 234.850000 87.530000 234.920000 ;
    END
  END key[85]
  PIN key[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 86.700000 234.850000 86.770000 234.920000 ;
    END
  END key[84]
  PIN key[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 85.940000 234.850000 86.010000 234.920000 ;
    END
  END key[83]
  PIN key[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 85.180000 234.850000 85.250000 234.920000 ;
    END
  END key[82]
  PIN key[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 84.420000 234.850000 84.490000 234.920000 ;
    END
  END key[81]
  PIN key[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 83.660000 234.850000 83.730000 234.920000 ;
    END
  END key[80]
  PIN key[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 82.900000 234.850000 82.970000 234.920000 ;
    END
  END key[79]
  PIN key[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 82.140000 234.850000 82.210000 234.920000 ;
    END
  END key[78]
  PIN key[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 81.380000 234.850000 81.450000 234.920000 ;
    END
  END key[77]
  PIN key[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 80.620000 234.850000 80.690000 234.920000 ;
    END
  END key[76]
  PIN key[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 79.860000 234.850000 79.930000 234.920000 ;
    END
  END key[75]
  PIN key[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 79.100000 234.850000 79.170000 234.920000 ;
    END
  END key[74]
  PIN key[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 78.340000 234.850000 78.410000 234.920000 ;
    END
  END key[73]
  PIN key[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 77.580000 234.850000 77.650000 234.920000 ;
    END
  END key[72]
  PIN key[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 76.820000 234.850000 76.890000 234.920000 ;
    END
  END key[71]
  PIN key[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 76.060000 234.850000 76.130000 234.920000 ;
    END
  END key[70]
  PIN key[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 75.300000 234.850000 75.370000 234.920000 ;
    END
  END key[69]
  PIN key[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 74.540000 234.850000 74.610000 234.920000 ;
    END
  END key[68]
  PIN key[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 73.780000 234.850000 73.850000 234.920000 ;
    END
  END key[67]
  PIN key[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 73.020000 234.850000 73.090000 234.920000 ;
    END
  END key[66]
  PIN key[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 72.260000 234.850000 72.330000 234.920000 ;
    END
  END key[65]
  PIN key[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 71.500000 234.850000 71.570000 234.920000 ;
    END
  END key[64]
  PIN key[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 70.740000 234.850000 70.810000 234.920000 ;
    END
  END key[63]
  PIN key[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 69.980000 234.850000 70.050000 234.920000 ;
    END
  END key[62]
  PIN key[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 69.220000 234.850000 69.290000 234.920000 ;
    END
  END key[61]
  PIN key[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 68.460000 234.850000 68.530000 234.920000 ;
    END
  END key[60]
  PIN key[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 67.700000 234.850000 67.770000 234.920000 ;
    END
  END key[59]
  PIN key[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 66.940000 234.850000 67.010000 234.920000 ;
    END
  END key[58]
  PIN key[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 66.180000 234.850000 66.250000 234.920000 ;
    END
  END key[57]
  PIN key[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 65.420000 234.850000 65.490000 234.920000 ;
    END
  END key[56]
  PIN key[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 64.660000 234.850000 64.730000 234.920000 ;
    END
  END key[55]
  PIN key[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 63.900000 234.850000 63.970000 234.920000 ;
    END
  END key[54]
  PIN key[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 63.140000 234.850000 63.210000 234.920000 ;
    END
  END key[53]
  PIN key[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 62.380000 234.850000 62.450000 234.920000 ;
    END
  END key[52]
  PIN key[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 61.620000 234.850000 61.690000 234.920000 ;
    END
  END key[51]
  PIN key[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 60.860000 234.850000 60.930000 234.920000 ;
    END
  END key[50]
  PIN key[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 60.100000 234.850000 60.170000 234.920000 ;
    END
  END key[49]
  PIN key[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 59.340000 234.850000 59.410000 234.920000 ;
    END
  END key[48]
  PIN key[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 58.580000 234.850000 58.650000 234.920000 ;
    END
  END key[47]
  PIN key[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 57.820000 234.850000 57.890000 234.920000 ;
    END
  END key[46]
  PIN key[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 57.060000 234.850000 57.130000 234.920000 ;
    END
  END key[45]
  PIN key[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 56.300000 234.850000 56.370000 234.920000 ;
    END
  END key[44]
  PIN key[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 55.540000 234.850000 55.610000 234.920000 ;
    END
  END key[43]
  PIN key[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 54.780000 234.850000 54.850000 234.920000 ;
    END
  END key[42]
  PIN key[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 54.020000 234.850000 54.090000 234.920000 ;
    END
  END key[41]
  PIN key[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 53.260000 234.850000 53.330000 234.920000 ;
    END
  END key[40]
  PIN key[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 52.500000 234.850000 52.570000 234.920000 ;
    END
  END key[39]
  PIN key[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 51.740000 234.850000 51.810000 234.920000 ;
    END
  END key[38]
  PIN key[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 50.980000 234.850000 51.050000 234.920000 ;
    END
  END key[37]
  PIN key[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 50.220000 234.850000 50.290000 234.920000 ;
    END
  END key[36]
  PIN key[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 49.460000 234.850000 49.530000 234.920000 ;
    END
  END key[35]
  PIN key[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 48.700000 234.850000 48.770000 234.920000 ;
    END
  END key[34]
  PIN key[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 47.940000 234.850000 48.010000 234.920000 ;
    END
  END key[33]
  PIN key[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 47.180000 234.850000 47.250000 234.920000 ;
    END
  END key[32]
  PIN key[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 46.420000 234.850000 46.490000 234.920000 ;
    END
  END key[31]
  PIN key[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 45.660000 234.850000 45.730000 234.920000 ;
    END
  END key[30]
  PIN key[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 44.900000 234.850000 44.970000 234.920000 ;
    END
  END key[29]
  PIN key[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 44.140000 234.850000 44.210000 234.920000 ;
    END
  END key[28]
  PIN key[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 43.380000 234.850000 43.450000 234.920000 ;
    END
  END key[27]
  PIN key[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 42.620000 234.850000 42.690000 234.920000 ;
    END
  END key[26]
  PIN key[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 41.860000 234.850000 41.930000 234.920000 ;
    END
  END key[25]
  PIN key[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 41.100000 234.850000 41.170000 234.920000 ;
    END
  END key[24]
  PIN key[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 40.340000 234.850000 40.410000 234.920000 ;
    END
  END key[23]
  PIN key[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 39.580000 234.850000 39.650000 234.920000 ;
    END
  END key[22]
  PIN key[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 38.820000 234.850000 38.890000 234.920000 ;
    END
  END key[21]
  PIN key[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 38.060000 234.850000 38.130000 234.920000 ;
    END
  END key[20]
  PIN key[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 37.300000 234.850000 37.370000 234.920000 ;
    END
  END key[19]
  PIN key[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 36.540000 234.850000 36.610000 234.920000 ;
    END
  END key[18]
  PIN key[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 35.780000 234.850000 35.850000 234.920000 ;
    END
  END key[17]
  PIN key[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 35.020000 234.850000 35.090000 234.920000 ;
    END
  END key[16]
  PIN key[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 34.260000 234.850000 34.330000 234.920000 ;
    END
  END key[15]
  PIN key[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 33.500000 234.850000 33.570000 234.920000 ;
    END
  END key[14]
  PIN key[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 32.740000 234.850000 32.810000 234.920000 ;
    END
  END key[13]
  PIN key[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 31.980000 234.850000 32.050000 234.920000 ;
    END
  END key[12]
  PIN key[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 31.220000 234.850000 31.290000 234.920000 ;
    END
  END key[11]
  PIN key[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 30.460000 234.850000 30.530000 234.920000 ;
    END
  END key[10]
  PIN key[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 29.700000 234.850000 29.770000 234.920000 ;
    END
  END key[9]
  PIN key[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 28.940000 234.850000 29.010000 234.920000 ;
    END
  END key[8]
  PIN key[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 28.180000 234.850000 28.250000 234.920000 ;
    END
  END key[7]
  PIN key[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 27.420000 234.850000 27.490000 234.920000 ;
    END
  END key[6]
  PIN key[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 26.660000 234.850000 26.730000 234.920000 ;
    END
  END key[5]
  PIN key[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 25.900000 234.850000 25.970000 234.920000 ;
    END
  END key[4]
  PIN key[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 25.140000 234.850000 25.210000 234.920000 ;
    END
  END key[3]
  PIN key[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 24.380000 234.850000 24.450000 234.920000 ;
    END
  END key[2]
  PIN key[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 23.620000 234.850000 23.690000 234.920000 ;
    END
  END key[1]
  PIN key[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 22.860000 234.850000 22.930000 234.920000 ;
    END
  END key[0]
  PIN plain[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 216.660000 234.850000 216.730000 234.920000 ;
    END
  END plain[127]
  PIN plain[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 215.900000 234.850000 215.970000 234.920000 ;
    END
  END plain[126]
  PIN plain[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 215.140000 234.850000 215.210000 234.920000 ;
    END
  END plain[125]
  PIN plain[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 214.380000 234.850000 214.450000 234.920000 ;
    END
  END plain[124]
  PIN plain[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 213.620000 234.850000 213.690000 234.920000 ;
    END
  END plain[123]
  PIN plain[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 212.860000 234.850000 212.930000 234.920000 ;
    END
  END plain[122]
  PIN plain[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 212.100000 234.850000 212.170000 234.920000 ;
    END
  END plain[121]
  PIN plain[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 211.340000 234.850000 211.410000 234.920000 ;
    END
  END plain[120]
  PIN plain[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 210.580000 234.850000 210.650000 234.920000 ;
    END
  END plain[119]
  PIN plain[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 209.820000 234.850000 209.890000 234.920000 ;
    END
  END plain[118]
  PIN plain[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 209.060000 234.850000 209.130000 234.920000 ;
    END
  END plain[117]
  PIN plain[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 208.300000 234.850000 208.370000 234.920000 ;
    END
  END plain[116]
  PIN plain[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 207.540000 234.850000 207.610000 234.920000 ;
    END
  END plain[115]
  PIN plain[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 206.780000 234.850000 206.850000 234.920000 ;
    END
  END plain[114]
  PIN plain[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 206.020000 234.850000 206.090000 234.920000 ;
    END
  END plain[113]
  PIN plain[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 205.260000 234.850000 205.330000 234.920000 ;
    END
  END plain[112]
  PIN plain[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 204.500000 234.850000 204.570000 234.920000 ;
    END
  END plain[111]
  PIN plain[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 203.740000 234.850000 203.810000 234.920000 ;
    END
  END plain[110]
  PIN plain[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 202.980000 234.850000 203.050000 234.920000 ;
    END
  END plain[109]
  PIN plain[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 202.220000 234.850000 202.290000 234.920000 ;
    END
  END plain[108]
  PIN plain[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 201.460000 234.850000 201.530000 234.920000 ;
    END
  END plain[107]
  PIN plain[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 200.700000 234.850000 200.770000 234.920000 ;
    END
  END plain[106]
  PIN plain[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 199.940000 234.850000 200.010000 234.920000 ;
    END
  END plain[105]
  PIN plain[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 199.180000 234.850000 199.250000 234.920000 ;
    END
  END plain[104]
  PIN plain[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 198.420000 234.850000 198.490000 234.920000 ;
    END
  END plain[103]
  PIN plain[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 197.660000 234.850000 197.730000 234.920000 ;
    END
  END plain[102]
  PIN plain[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 196.900000 234.850000 196.970000 234.920000 ;
    END
  END plain[101]
  PIN plain[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 196.140000 234.850000 196.210000 234.920000 ;
    END
  END plain[100]
  PIN plain[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 195.380000 234.850000 195.450000 234.920000 ;
    END
  END plain[99]
  PIN plain[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 194.620000 234.850000 194.690000 234.920000 ;
    END
  END plain[98]
  PIN plain[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 193.860000 234.850000 193.930000 234.920000 ;
    END
  END plain[97]
  PIN plain[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 193.100000 234.850000 193.170000 234.920000 ;
    END
  END plain[96]
  PIN plain[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 192.340000 234.850000 192.410000 234.920000 ;
    END
  END plain[95]
  PIN plain[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 191.580000 234.850000 191.650000 234.920000 ;
    END
  END plain[94]
  PIN plain[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 190.820000 234.850000 190.890000 234.920000 ;
    END
  END plain[93]
  PIN plain[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 190.060000 234.850000 190.130000 234.920000 ;
    END
  END plain[92]
  PIN plain[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 189.300000 234.850000 189.370000 234.920000 ;
    END
  END plain[91]
  PIN plain[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 188.540000 234.850000 188.610000 234.920000 ;
    END
  END plain[90]
  PIN plain[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 187.780000 234.850000 187.850000 234.920000 ;
    END
  END plain[89]
  PIN plain[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 187.020000 234.850000 187.090000 234.920000 ;
    END
  END plain[88]
  PIN plain[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 186.260000 234.850000 186.330000 234.920000 ;
    END
  END plain[87]
  PIN plain[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 185.500000 234.850000 185.570000 234.920000 ;
    END
  END plain[86]
  PIN plain[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 184.740000 234.850000 184.810000 234.920000 ;
    END
  END plain[85]
  PIN plain[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 183.980000 234.850000 184.050000 234.920000 ;
    END
  END plain[84]
  PIN plain[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 183.220000 234.850000 183.290000 234.920000 ;
    END
  END plain[83]
  PIN plain[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 182.460000 234.850000 182.530000 234.920000 ;
    END
  END plain[82]
  PIN plain[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 181.700000 234.850000 181.770000 234.920000 ;
    END
  END plain[81]
  PIN plain[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 180.940000 234.850000 181.010000 234.920000 ;
    END
  END plain[80]
  PIN plain[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 180.180000 234.850000 180.250000 234.920000 ;
    END
  END plain[79]
  PIN plain[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 179.420000 234.850000 179.490000 234.920000 ;
    END
  END plain[78]
  PIN plain[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 178.660000 234.850000 178.730000 234.920000 ;
    END
  END plain[77]
  PIN plain[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 177.900000 234.850000 177.970000 234.920000 ;
    END
  END plain[76]
  PIN plain[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 177.140000 234.850000 177.210000 234.920000 ;
    END
  END plain[75]
  PIN plain[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 176.380000 234.850000 176.450000 234.920000 ;
    END
  END plain[74]
  PIN plain[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 175.620000 234.850000 175.690000 234.920000 ;
    END
  END plain[73]
  PIN plain[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 174.860000 234.850000 174.930000 234.920000 ;
    END
  END plain[72]
  PIN plain[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 174.100000 234.850000 174.170000 234.920000 ;
    END
  END plain[71]
  PIN plain[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 173.340000 234.850000 173.410000 234.920000 ;
    END
  END plain[70]
  PIN plain[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 172.580000 234.850000 172.650000 234.920000 ;
    END
  END plain[69]
  PIN plain[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 171.820000 234.850000 171.890000 234.920000 ;
    END
  END plain[68]
  PIN plain[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 171.060000 234.850000 171.130000 234.920000 ;
    END
  END plain[67]
  PIN plain[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 170.300000 234.850000 170.370000 234.920000 ;
    END
  END plain[66]
  PIN plain[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 169.540000 234.850000 169.610000 234.920000 ;
    END
  END plain[65]
  PIN plain[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 168.780000 234.850000 168.850000 234.920000 ;
    END
  END plain[64]
  PIN plain[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 168.020000 234.850000 168.090000 234.920000 ;
    END
  END plain[63]
  PIN plain[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 167.260000 234.850000 167.330000 234.920000 ;
    END
  END plain[62]
  PIN plain[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 166.500000 234.850000 166.570000 234.920000 ;
    END
  END plain[61]
  PIN plain[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 165.740000 234.850000 165.810000 234.920000 ;
    END
  END plain[60]
  PIN plain[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 164.980000 234.850000 165.050000 234.920000 ;
    END
  END plain[59]
  PIN plain[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 164.220000 234.850000 164.290000 234.920000 ;
    END
  END plain[58]
  PIN plain[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 163.460000 234.850000 163.530000 234.920000 ;
    END
  END plain[57]
  PIN plain[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 162.700000 234.850000 162.770000 234.920000 ;
    END
  END plain[56]
  PIN plain[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 161.940000 234.850000 162.010000 234.920000 ;
    END
  END plain[55]
  PIN plain[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 161.180000 234.850000 161.250000 234.920000 ;
    END
  END plain[54]
  PIN plain[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 160.420000 234.850000 160.490000 234.920000 ;
    END
  END plain[53]
  PIN plain[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 159.660000 234.850000 159.730000 234.920000 ;
    END
  END plain[52]
  PIN plain[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 158.900000 234.850000 158.970000 234.920000 ;
    END
  END plain[51]
  PIN plain[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 158.140000 234.850000 158.210000 234.920000 ;
    END
  END plain[50]
  PIN plain[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 157.380000 234.850000 157.450000 234.920000 ;
    END
  END plain[49]
  PIN plain[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 156.620000 234.850000 156.690000 234.920000 ;
    END
  END plain[48]
  PIN plain[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 155.860000 234.850000 155.930000 234.920000 ;
    END
  END plain[47]
  PIN plain[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 155.100000 234.850000 155.170000 234.920000 ;
    END
  END plain[46]
  PIN plain[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 154.340000 234.850000 154.410000 234.920000 ;
    END
  END plain[45]
  PIN plain[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 153.580000 234.850000 153.650000 234.920000 ;
    END
  END plain[44]
  PIN plain[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 152.820000 234.850000 152.890000 234.920000 ;
    END
  END plain[43]
  PIN plain[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 152.060000 234.850000 152.130000 234.920000 ;
    END
  END plain[42]
  PIN plain[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 151.300000 234.850000 151.370000 234.920000 ;
    END
  END plain[41]
  PIN plain[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 150.540000 234.850000 150.610000 234.920000 ;
    END
  END plain[40]
  PIN plain[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 149.780000 234.850000 149.850000 234.920000 ;
    END
  END plain[39]
  PIN plain[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 149.020000 234.850000 149.090000 234.920000 ;
    END
  END plain[38]
  PIN plain[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 148.260000 234.850000 148.330000 234.920000 ;
    END
  END plain[37]
  PIN plain[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 147.500000 234.850000 147.570000 234.920000 ;
    END
  END plain[36]
  PIN plain[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 146.740000 234.850000 146.810000 234.920000 ;
    END
  END plain[35]
  PIN plain[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 145.980000 234.850000 146.050000 234.920000 ;
    END
  END plain[34]
  PIN plain[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 145.220000 234.850000 145.290000 234.920000 ;
    END
  END plain[33]
  PIN plain[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 144.460000 234.850000 144.530000 234.920000 ;
    END
  END plain[32]
  PIN plain[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 143.700000 234.850000 143.770000 234.920000 ;
    END
  END plain[31]
  PIN plain[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 142.940000 234.850000 143.010000 234.920000 ;
    END
  END plain[30]
  PIN plain[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 142.180000 234.850000 142.250000 234.920000 ;
    END
  END plain[29]
  PIN plain[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 141.420000 234.850000 141.490000 234.920000 ;
    END
  END plain[28]
  PIN plain[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 140.660000 234.850000 140.730000 234.920000 ;
    END
  END plain[27]
  PIN plain[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 139.900000 234.850000 139.970000 234.920000 ;
    END
  END plain[26]
  PIN plain[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 139.140000 234.850000 139.210000 234.920000 ;
    END
  END plain[25]
  PIN plain[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 138.380000 234.850000 138.450000 234.920000 ;
    END
  END plain[24]
  PIN plain[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 137.620000 234.850000 137.690000 234.920000 ;
    END
  END plain[23]
  PIN plain[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 136.860000 234.850000 136.930000 234.920000 ;
    END
  END plain[22]
  PIN plain[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 136.100000 234.850000 136.170000 234.920000 ;
    END
  END plain[21]
  PIN plain[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 135.340000 234.850000 135.410000 234.920000 ;
    END
  END plain[20]
  PIN plain[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 134.580000 234.850000 134.650000 234.920000 ;
    END
  END plain[19]
  PIN plain[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 133.820000 234.850000 133.890000 234.920000 ;
    END
  END plain[18]
  PIN plain[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 133.060000 234.850000 133.130000 234.920000 ;
    END
  END plain[17]
  PIN plain[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 132.300000 234.850000 132.370000 234.920000 ;
    END
  END plain[16]
  PIN plain[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 131.540000 234.850000 131.610000 234.920000 ;
    END
  END plain[15]
  PIN plain[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 130.780000 234.850000 130.850000 234.920000 ;
    END
  END plain[14]
  PIN plain[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 130.020000 234.850000 130.090000 234.920000 ;
    END
  END plain[13]
  PIN plain[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 129.260000 234.850000 129.330000 234.920000 ;
    END
  END plain[12]
  PIN plain[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 128.500000 234.850000 128.570000 234.920000 ;
    END
  END plain[11]
  PIN plain[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 127.740000 234.850000 127.810000 234.920000 ;
    END
  END plain[10]
  PIN plain[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 126.980000 234.850000 127.050000 234.920000 ;
    END
  END plain[9]
  PIN plain[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 126.220000 234.850000 126.290000 234.920000 ;
    END
  END plain[8]
  PIN plain[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 125.460000 234.850000 125.530000 234.920000 ;
    END
  END plain[7]
  PIN plain[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 124.700000 234.850000 124.770000 234.920000 ;
    END
  END plain[6]
  PIN plain[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 123.940000 234.850000 124.010000 234.920000 ;
    END
  END plain[5]
  PIN plain[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 123.180000 234.850000 123.250000 234.920000 ;
    END
  END plain[4]
  PIN plain[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 122.420000 234.850000 122.490000 234.920000 ;
    END
  END plain[3]
  PIN plain[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 121.660000 234.850000 121.730000 234.920000 ;
    END
  END plain[2]
  PIN plain[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 120.900000 234.850000 120.970000 234.920000 ;
    END
  END plain[1]
  PIN plain[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 120.140000 234.850000 120.210000 234.920000 ;
    END
  END plain[0]
  PIN ready
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 228.060000 0.000000 228.130000 0.070000 ;
    END
  END ready
  PIN cipher[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 9.180000 0.000000 9.250000 0.070000 ;
    END
  END cipher[127]
  PIN cipher[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 10.890000 0.000000 10.960000 0.070000 ;
    END
  END cipher[126]
  PIN cipher[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 12.600000 0.000000 12.670000 0.070000 ;
    END
  END cipher[125]
  PIN cipher[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 14.310000 0.000000 14.380000 0.070000 ;
    END
  END cipher[124]
  PIN cipher[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 16.020000 0.000000 16.090000 0.070000 ;
    END
  END cipher[123]
  PIN cipher[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 17.730000 0.000000 17.800000 0.070000 ;
    END
  END cipher[122]
  PIN cipher[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 19.440000 0.000000 19.510000 0.070000 ;
    END
  END cipher[121]
  PIN cipher[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 21.150000 0.000000 21.220000 0.070000 ;
    END
  END cipher[120]
  PIN cipher[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 22.860000 0.000000 22.930000 0.070000 ;
    END
  END cipher[119]
  PIN cipher[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 24.570000 0.000000 24.640000 0.070000 ;
    END
  END cipher[118]
  PIN cipher[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 26.280000 0.000000 26.350000 0.070000 ;
    END
  END cipher[117]
  PIN cipher[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 27.990000 0.000000 28.060000 0.070000 ;
    END
  END cipher[116]
  PIN cipher[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 29.700000 0.000000 29.770000 0.070000 ;
    END
  END cipher[115]
  PIN cipher[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 31.410000 0.000000 31.480000 0.070000 ;
    END
  END cipher[114]
  PIN cipher[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 33.120000 0.000000 33.190000 0.070000 ;
    END
  END cipher[113]
  PIN cipher[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 34.830000 0.000000 34.900000 0.070000 ;
    END
  END cipher[112]
  PIN cipher[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 36.540000 0.000000 36.610000 0.070000 ;
    END
  END cipher[111]
  PIN cipher[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 38.250000 0.000000 38.320000 0.070000 ;
    END
  END cipher[110]
  PIN cipher[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 39.960000 0.000000 40.030000 0.070000 ;
    END
  END cipher[109]
  PIN cipher[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 41.670000 0.000000 41.740000 0.070000 ;
    END
  END cipher[108]
  PIN cipher[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 43.380000 0.000000 43.450000 0.070000 ;
    END
  END cipher[107]
  PIN cipher[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 45.090000 0.000000 45.160000 0.070000 ;
    END
  END cipher[106]
  PIN cipher[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 46.800000 0.000000 46.870000 0.070000 ;
    END
  END cipher[105]
  PIN cipher[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 48.510000 0.000000 48.580000 0.070000 ;
    END
  END cipher[104]
  PIN cipher[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 50.220000 0.000000 50.290000 0.070000 ;
    END
  END cipher[103]
  PIN cipher[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 51.930000 0.000000 52.000000 0.070000 ;
    END
  END cipher[102]
  PIN cipher[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 53.640000 0.000000 53.710000 0.070000 ;
    END
  END cipher[101]
  PIN cipher[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 55.350000 0.000000 55.420000 0.070000 ;
    END
  END cipher[100]
  PIN cipher[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 57.060000 0.000000 57.130000 0.070000 ;
    END
  END cipher[99]
  PIN cipher[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 58.770000 0.000000 58.840000 0.070000 ;
    END
  END cipher[98]
  PIN cipher[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 60.480000 0.000000 60.550000 0.070000 ;
    END
  END cipher[97]
  PIN cipher[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 62.190000 0.000000 62.260000 0.070000 ;
    END
  END cipher[96]
  PIN cipher[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 63.900000 0.000000 63.970000 0.070000 ;
    END
  END cipher[95]
  PIN cipher[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 65.610000 0.000000 65.680000 0.070000 ;
    END
  END cipher[94]
  PIN cipher[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 67.320000 0.000000 67.390000 0.070000 ;
    END
  END cipher[93]
  PIN cipher[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 69.030000 0.000000 69.100000 0.070000 ;
    END
  END cipher[92]
  PIN cipher[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 70.740000 0.000000 70.810000 0.070000 ;
    END
  END cipher[91]
  PIN cipher[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 72.450000 0.000000 72.520000 0.070000 ;
    END
  END cipher[90]
  PIN cipher[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 74.160000 0.000000 74.230000 0.070000 ;
    END
  END cipher[89]
  PIN cipher[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 75.870000 0.000000 75.940000 0.070000 ;
    END
  END cipher[88]
  PIN cipher[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 77.580000 0.000000 77.650000 0.070000 ;
    END
  END cipher[87]
  PIN cipher[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 79.290000 0.000000 79.360000 0.070000 ;
    END
  END cipher[86]
  PIN cipher[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 81.000000 0.000000 81.070000 0.070000 ;
    END
  END cipher[85]
  PIN cipher[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 82.710000 0.000000 82.780000 0.070000 ;
    END
  END cipher[84]
  PIN cipher[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 84.420000 0.000000 84.490000 0.070000 ;
    END
  END cipher[83]
  PIN cipher[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 86.130000 0.000000 86.200000 0.070000 ;
    END
  END cipher[82]
  PIN cipher[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 87.840000 0.000000 87.910000 0.070000 ;
    END
  END cipher[81]
  PIN cipher[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 89.550000 0.000000 89.620000 0.070000 ;
    END
  END cipher[80]
  PIN cipher[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 91.260000 0.000000 91.330000 0.070000 ;
    END
  END cipher[79]
  PIN cipher[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 92.970000 0.000000 93.040000 0.070000 ;
    END
  END cipher[78]
  PIN cipher[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 94.680000 0.000000 94.750000 0.070000 ;
    END
  END cipher[77]
  PIN cipher[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 96.390000 0.000000 96.460000 0.070000 ;
    END
  END cipher[76]
  PIN cipher[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 98.100000 0.000000 98.170000 0.070000 ;
    END
  END cipher[75]
  PIN cipher[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 99.810000 0.000000 99.880000 0.070000 ;
    END
  END cipher[74]
  PIN cipher[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 101.520000 0.000000 101.590000 0.070000 ;
    END
  END cipher[73]
  PIN cipher[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 103.230000 0.000000 103.300000 0.070000 ;
    END
  END cipher[72]
  PIN cipher[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 104.940000 0.000000 105.010000 0.070000 ;
    END
  END cipher[71]
  PIN cipher[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 106.650000 0.000000 106.720000 0.070000 ;
    END
  END cipher[70]
  PIN cipher[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 108.360000 0.000000 108.430000 0.070000 ;
    END
  END cipher[69]
  PIN cipher[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 110.070000 0.000000 110.140000 0.070000 ;
    END
  END cipher[68]
  PIN cipher[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 111.780000 0.000000 111.850000 0.070000 ;
    END
  END cipher[67]
  PIN cipher[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 113.490000 0.000000 113.560000 0.070000 ;
    END
  END cipher[66]
  PIN cipher[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 115.200000 0.000000 115.270000 0.070000 ;
    END
  END cipher[65]
  PIN cipher[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 116.910000 0.000000 116.980000 0.070000 ;
    END
  END cipher[64]
  PIN cipher[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 118.620000 0.000000 118.690000 0.070000 ;
    END
  END cipher[63]
  PIN cipher[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 120.330000 0.000000 120.400000 0.070000 ;
    END
  END cipher[62]
  PIN cipher[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 122.040000 0.000000 122.110000 0.070000 ;
    END
  END cipher[61]
  PIN cipher[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 123.750000 0.000000 123.820000 0.070000 ;
    END
  END cipher[60]
  PIN cipher[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 125.460000 0.000000 125.530000 0.070000 ;
    END
  END cipher[59]
  PIN cipher[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 127.170000 0.000000 127.240000 0.070000 ;
    END
  END cipher[58]
  PIN cipher[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 128.880000 0.000000 128.950000 0.070000 ;
    END
  END cipher[57]
  PIN cipher[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 130.590000 0.000000 130.660000 0.070000 ;
    END
  END cipher[56]
  PIN cipher[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 132.300000 0.000000 132.370000 0.070000 ;
    END
  END cipher[55]
  PIN cipher[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 134.010000 0.000000 134.080000 0.070000 ;
    END
  END cipher[54]
  PIN cipher[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 135.720000 0.000000 135.790000 0.070000 ;
    END
  END cipher[53]
  PIN cipher[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 137.430000 0.000000 137.500000 0.070000 ;
    END
  END cipher[52]
  PIN cipher[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 139.140000 0.000000 139.210000 0.070000 ;
    END
  END cipher[51]
  PIN cipher[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 140.850000 0.000000 140.920000 0.070000 ;
    END
  END cipher[50]
  PIN cipher[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 142.560000 0.000000 142.630000 0.070000 ;
    END
  END cipher[49]
  PIN cipher[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 144.270000 0.000000 144.340000 0.070000 ;
    END
  END cipher[48]
  PIN cipher[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 145.980000 0.000000 146.050000 0.070000 ;
    END
  END cipher[47]
  PIN cipher[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 147.690000 0.000000 147.760000 0.070000 ;
    END
  END cipher[46]
  PIN cipher[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 149.400000 0.000000 149.470000 0.070000 ;
    END
  END cipher[45]
  PIN cipher[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 151.110000 0.000000 151.180000 0.070000 ;
    END
  END cipher[44]
  PIN cipher[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 152.820000 0.000000 152.890000 0.070000 ;
    END
  END cipher[43]
  PIN cipher[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 154.530000 0.000000 154.600000 0.070000 ;
    END
  END cipher[42]
  PIN cipher[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 156.240000 0.000000 156.310000 0.070000 ;
    END
  END cipher[41]
  PIN cipher[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 157.950000 0.000000 158.020000 0.070000 ;
    END
  END cipher[40]
  PIN cipher[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 159.660000 0.000000 159.730000 0.070000 ;
    END
  END cipher[39]
  PIN cipher[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 161.370000 0.000000 161.440000 0.070000 ;
    END
  END cipher[38]
  PIN cipher[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 163.080000 0.000000 163.150000 0.070000 ;
    END
  END cipher[37]
  PIN cipher[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 164.790000 0.000000 164.860000 0.070000 ;
    END
  END cipher[36]
  PIN cipher[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 166.500000 0.000000 166.570000 0.070000 ;
    END
  END cipher[35]
  PIN cipher[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 168.210000 0.000000 168.280000 0.070000 ;
    END
  END cipher[34]
  PIN cipher[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 169.920000 0.000000 169.990000 0.070000 ;
    END
  END cipher[33]
  PIN cipher[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 171.630000 0.000000 171.700000 0.070000 ;
    END
  END cipher[32]
  PIN cipher[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 173.340000 0.000000 173.410000 0.070000 ;
    END
  END cipher[31]
  PIN cipher[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 175.050000 0.000000 175.120000 0.070000 ;
    END
  END cipher[30]
  PIN cipher[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 176.760000 0.000000 176.830000 0.070000 ;
    END
  END cipher[29]
  PIN cipher[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 178.470000 0.000000 178.540000 0.070000 ;
    END
  END cipher[28]
  PIN cipher[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 180.180000 0.000000 180.250000 0.070000 ;
    END
  END cipher[27]
  PIN cipher[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 181.890000 0.000000 181.960000 0.070000 ;
    END
  END cipher[26]
  PIN cipher[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 183.600000 0.000000 183.670000 0.070000 ;
    END
  END cipher[25]
  PIN cipher[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 185.310000 0.000000 185.380000 0.070000 ;
    END
  END cipher[24]
  PIN cipher[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 187.020000 0.000000 187.090000 0.070000 ;
    END
  END cipher[23]
  PIN cipher[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 188.730000 0.000000 188.800000 0.070000 ;
    END
  END cipher[22]
  PIN cipher[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 190.440000 0.000000 190.510000 0.070000 ;
    END
  END cipher[21]
  PIN cipher[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 192.150000 0.000000 192.220000 0.070000 ;
    END
  END cipher[20]
  PIN cipher[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 193.860000 0.000000 193.930000 0.070000 ;
    END
  END cipher[19]
  PIN cipher[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 195.570000 0.000000 195.640000 0.070000 ;
    END
  END cipher[18]
  PIN cipher[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 197.280000 0.000000 197.350000 0.070000 ;
    END
  END cipher[17]
  PIN cipher[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 198.990000 0.000000 199.060000 0.070000 ;
    END
  END cipher[16]
  PIN cipher[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 200.700000 0.000000 200.770000 0.070000 ;
    END
  END cipher[15]
  PIN cipher[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 202.410000 0.000000 202.480000 0.070000 ;
    END
  END cipher[14]
  PIN cipher[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 204.120000 0.000000 204.190000 0.070000 ;
    END
  END cipher[13]
  PIN cipher[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 205.830000 0.000000 205.900000 0.070000 ;
    END
  END cipher[12]
  PIN cipher[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 207.540000 0.000000 207.610000 0.070000 ;
    END
  END cipher[11]
  PIN cipher[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 209.250000 0.000000 209.320000 0.070000 ;
    END
  END cipher[10]
  PIN cipher[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 210.960000 0.000000 211.030000 0.070000 ;
    END
  END cipher[9]
  PIN cipher[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 212.670000 0.000000 212.740000 0.070000 ;
    END
  END cipher[8]
  PIN cipher[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 214.380000 0.000000 214.450000 0.070000 ;
    END
  END cipher[7]
  PIN cipher[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 216.090000 0.000000 216.160000 0.070000 ;
    END
  END cipher[6]
  PIN cipher[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 217.800000 0.000000 217.870000 0.070000 ;
    END
  END cipher[5]
  PIN cipher[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 219.510000 0.000000 219.580000 0.070000 ;
    END
  END cipher[4]
  PIN cipher[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 221.220000 0.000000 221.290000 0.070000 ;
    END
  END cipher[3]
  PIN cipher[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 222.930000 0.000000 223.000000 0.070000 ;
    END
  END cipher[2]
  PIN cipher[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 224.640000 0.000000 224.710000 0.070000 ;
    END
  END cipher[1]
  PIN cipher[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 226.350000 0.000000 226.420000 0.070000 ;
    END
  END cipher[0]
  OBS
    LAYER metal1 ;
      RECT 0.000000 0.000000 236.930000 234.920000 ;
    LAYER metal2 ;
      RECT 216.800000 234.780000 236.930000 234.920000 ;
      RECT 216.040000 234.780000 216.590000 234.920000 ;
      RECT 215.280000 234.780000 215.830000 234.920000 ;
      RECT 214.520000 234.780000 215.070000 234.920000 ;
      RECT 213.760000 234.780000 214.310000 234.920000 ;
      RECT 213.000000 234.780000 213.550000 234.920000 ;
      RECT 212.240000 234.780000 212.790000 234.920000 ;
      RECT 211.480000 234.780000 212.030000 234.920000 ;
      RECT 210.720000 234.780000 211.270000 234.920000 ;
      RECT 209.960000 234.780000 210.510000 234.920000 ;
      RECT 209.200000 234.780000 209.750000 234.920000 ;
      RECT 208.440000 234.780000 208.990000 234.920000 ;
      RECT 207.680000 234.780000 208.230000 234.920000 ;
      RECT 206.920000 234.780000 207.470000 234.920000 ;
      RECT 206.160000 234.780000 206.710000 234.920000 ;
      RECT 205.400000 234.780000 205.950000 234.920000 ;
      RECT 204.640000 234.780000 205.190000 234.920000 ;
      RECT 203.880000 234.780000 204.430000 234.920000 ;
      RECT 203.120000 234.780000 203.670000 234.920000 ;
      RECT 202.360000 234.780000 202.910000 234.920000 ;
      RECT 201.600000 234.780000 202.150000 234.920000 ;
      RECT 200.840000 234.780000 201.390000 234.920000 ;
      RECT 200.080000 234.780000 200.630000 234.920000 ;
      RECT 199.320000 234.780000 199.870000 234.920000 ;
      RECT 198.560000 234.780000 199.110000 234.920000 ;
      RECT 197.800000 234.780000 198.350000 234.920000 ;
      RECT 197.040000 234.780000 197.590000 234.920000 ;
      RECT 196.280000 234.780000 196.830000 234.920000 ;
      RECT 195.520000 234.780000 196.070000 234.920000 ;
      RECT 194.760000 234.780000 195.310000 234.920000 ;
      RECT 194.000000 234.780000 194.550000 234.920000 ;
      RECT 193.240000 234.780000 193.790000 234.920000 ;
      RECT 192.480000 234.780000 193.030000 234.920000 ;
      RECT 191.720000 234.780000 192.270000 234.920000 ;
      RECT 190.960000 234.780000 191.510000 234.920000 ;
      RECT 190.200000 234.780000 190.750000 234.920000 ;
      RECT 189.440000 234.780000 189.990000 234.920000 ;
      RECT 188.680000 234.780000 189.230000 234.920000 ;
      RECT 187.920000 234.780000 188.470000 234.920000 ;
      RECT 187.160000 234.780000 187.710000 234.920000 ;
      RECT 186.400000 234.780000 186.950000 234.920000 ;
      RECT 185.640000 234.780000 186.190000 234.920000 ;
      RECT 184.880000 234.780000 185.430000 234.920000 ;
      RECT 184.120000 234.780000 184.670000 234.920000 ;
      RECT 183.360000 234.780000 183.910000 234.920000 ;
      RECT 182.600000 234.780000 183.150000 234.920000 ;
      RECT 181.840000 234.780000 182.390000 234.920000 ;
      RECT 181.080000 234.780000 181.630000 234.920000 ;
      RECT 180.320000 234.780000 180.870000 234.920000 ;
      RECT 179.560000 234.780000 180.110000 234.920000 ;
      RECT 178.800000 234.780000 179.350000 234.920000 ;
      RECT 178.040000 234.780000 178.590000 234.920000 ;
      RECT 177.280000 234.780000 177.830000 234.920000 ;
      RECT 176.520000 234.780000 177.070000 234.920000 ;
      RECT 175.760000 234.780000 176.310000 234.920000 ;
      RECT 175.000000 234.780000 175.550000 234.920000 ;
      RECT 174.240000 234.780000 174.790000 234.920000 ;
      RECT 173.480000 234.780000 174.030000 234.920000 ;
      RECT 172.720000 234.780000 173.270000 234.920000 ;
      RECT 171.960000 234.780000 172.510000 234.920000 ;
      RECT 171.200000 234.780000 171.750000 234.920000 ;
      RECT 170.440000 234.780000 170.990000 234.920000 ;
      RECT 169.680000 234.780000 170.230000 234.920000 ;
      RECT 168.920000 234.780000 169.470000 234.920000 ;
      RECT 168.160000 234.780000 168.710000 234.920000 ;
      RECT 167.400000 234.780000 167.950000 234.920000 ;
      RECT 166.640000 234.780000 167.190000 234.920000 ;
      RECT 165.880000 234.780000 166.430000 234.920000 ;
      RECT 165.120000 234.780000 165.670000 234.920000 ;
      RECT 164.360000 234.780000 164.910000 234.920000 ;
      RECT 163.600000 234.780000 164.150000 234.920000 ;
      RECT 162.840000 234.780000 163.390000 234.920000 ;
      RECT 162.080000 234.780000 162.630000 234.920000 ;
      RECT 161.320000 234.780000 161.870000 234.920000 ;
      RECT 160.560000 234.780000 161.110000 234.920000 ;
      RECT 159.800000 234.780000 160.350000 234.920000 ;
      RECT 159.040000 234.780000 159.590000 234.920000 ;
      RECT 158.280000 234.780000 158.830000 234.920000 ;
      RECT 157.520000 234.780000 158.070000 234.920000 ;
      RECT 156.760000 234.780000 157.310000 234.920000 ;
      RECT 156.000000 234.780000 156.550000 234.920000 ;
      RECT 155.240000 234.780000 155.790000 234.920000 ;
      RECT 154.480000 234.780000 155.030000 234.920000 ;
      RECT 153.720000 234.780000 154.270000 234.920000 ;
      RECT 152.960000 234.780000 153.510000 234.920000 ;
      RECT 152.200000 234.780000 152.750000 234.920000 ;
      RECT 151.440000 234.780000 151.990000 234.920000 ;
      RECT 150.680000 234.780000 151.230000 234.920000 ;
      RECT 149.920000 234.780000 150.470000 234.920000 ;
      RECT 149.160000 234.780000 149.710000 234.920000 ;
      RECT 148.400000 234.780000 148.950000 234.920000 ;
      RECT 147.640000 234.780000 148.190000 234.920000 ;
      RECT 146.880000 234.780000 147.430000 234.920000 ;
      RECT 146.120000 234.780000 146.670000 234.920000 ;
      RECT 145.360000 234.780000 145.910000 234.920000 ;
      RECT 144.600000 234.780000 145.150000 234.920000 ;
      RECT 143.840000 234.780000 144.390000 234.920000 ;
      RECT 143.080000 234.780000 143.630000 234.920000 ;
      RECT 142.320000 234.780000 142.870000 234.920000 ;
      RECT 141.560000 234.780000 142.110000 234.920000 ;
      RECT 140.800000 234.780000 141.350000 234.920000 ;
      RECT 140.040000 234.780000 140.590000 234.920000 ;
      RECT 139.280000 234.780000 139.830000 234.920000 ;
      RECT 138.520000 234.780000 139.070000 234.920000 ;
      RECT 137.760000 234.780000 138.310000 234.920000 ;
      RECT 137.000000 234.780000 137.550000 234.920000 ;
      RECT 136.240000 234.780000 136.790000 234.920000 ;
      RECT 135.480000 234.780000 136.030000 234.920000 ;
      RECT 134.720000 234.780000 135.270000 234.920000 ;
      RECT 133.960000 234.780000 134.510000 234.920000 ;
      RECT 133.200000 234.780000 133.750000 234.920000 ;
      RECT 132.440000 234.780000 132.990000 234.920000 ;
      RECT 131.680000 234.780000 132.230000 234.920000 ;
      RECT 130.920000 234.780000 131.470000 234.920000 ;
      RECT 130.160000 234.780000 130.710000 234.920000 ;
      RECT 129.400000 234.780000 129.950000 234.920000 ;
      RECT 128.640000 234.780000 129.190000 234.920000 ;
      RECT 127.880000 234.780000 128.430000 234.920000 ;
      RECT 127.120000 234.780000 127.670000 234.920000 ;
      RECT 126.360000 234.780000 126.910000 234.920000 ;
      RECT 125.600000 234.780000 126.150000 234.920000 ;
      RECT 124.840000 234.780000 125.390000 234.920000 ;
      RECT 124.080000 234.780000 124.630000 234.920000 ;
      RECT 123.320000 234.780000 123.870000 234.920000 ;
      RECT 122.560000 234.780000 123.110000 234.920000 ;
      RECT 121.800000 234.780000 122.350000 234.920000 ;
      RECT 121.040000 234.780000 121.590000 234.920000 ;
      RECT 120.280000 234.780000 120.830000 234.920000 ;
      RECT 119.520000 234.780000 120.070000 234.920000 ;
      RECT 118.760000 234.780000 119.310000 234.920000 ;
      RECT 118.000000 234.780000 118.550000 234.920000 ;
      RECT 117.240000 234.780000 117.790000 234.920000 ;
      RECT 116.480000 234.780000 117.030000 234.920000 ;
      RECT 115.720000 234.780000 116.270000 234.920000 ;
      RECT 114.960000 234.780000 115.510000 234.920000 ;
      RECT 114.200000 234.780000 114.750000 234.920000 ;
      RECT 113.440000 234.780000 113.990000 234.920000 ;
      RECT 112.680000 234.780000 113.230000 234.920000 ;
      RECT 111.920000 234.780000 112.470000 234.920000 ;
      RECT 111.160000 234.780000 111.710000 234.920000 ;
      RECT 110.400000 234.780000 110.950000 234.920000 ;
      RECT 109.640000 234.780000 110.190000 234.920000 ;
      RECT 108.880000 234.780000 109.430000 234.920000 ;
      RECT 108.120000 234.780000 108.670000 234.920000 ;
      RECT 107.360000 234.780000 107.910000 234.920000 ;
      RECT 106.600000 234.780000 107.150000 234.920000 ;
      RECT 105.840000 234.780000 106.390000 234.920000 ;
      RECT 105.080000 234.780000 105.630000 234.920000 ;
      RECT 104.320000 234.780000 104.870000 234.920000 ;
      RECT 103.560000 234.780000 104.110000 234.920000 ;
      RECT 102.800000 234.780000 103.350000 234.920000 ;
      RECT 102.040000 234.780000 102.590000 234.920000 ;
      RECT 101.280000 234.780000 101.830000 234.920000 ;
      RECT 100.520000 234.780000 101.070000 234.920000 ;
      RECT 99.760000 234.780000 100.310000 234.920000 ;
      RECT 99.000000 234.780000 99.550000 234.920000 ;
      RECT 98.240000 234.780000 98.790000 234.920000 ;
      RECT 97.480000 234.780000 98.030000 234.920000 ;
      RECT 96.720000 234.780000 97.270000 234.920000 ;
      RECT 95.960000 234.780000 96.510000 234.920000 ;
      RECT 95.200000 234.780000 95.750000 234.920000 ;
      RECT 94.440000 234.780000 94.990000 234.920000 ;
      RECT 93.680000 234.780000 94.230000 234.920000 ;
      RECT 92.920000 234.780000 93.470000 234.920000 ;
      RECT 92.160000 234.780000 92.710000 234.920000 ;
      RECT 91.400000 234.780000 91.950000 234.920000 ;
      RECT 90.640000 234.780000 91.190000 234.920000 ;
      RECT 89.880000 234.780000 90.430000 234.920000 ;
      RECT 89.120000 234.780000 89.670000 234.920000 ;
      RECT 88.360000 234.780000 88.910000 234.920000 ;
      RECT 87.600000 234.780000 88.150000 234.920000 ;
      RECT 86.840000 234.780000 87.390000 234.920000 ;
      RECT 86.080000 234.780000 86.630000 234.920000 ;
      RECT 85.320000 234.780000 85.870000 234.920000 ;
      RECT 84.560000 234.780000 85.110000 234.920000 ;
      RECT 83.800000 234.780000 84.350000 234.920000 ;
      RECT 83.040000 234.780000 83.590000 234.920000 ;
      RECT 82.280000 234.780000 82.830000 234.920000 ;
      RECT 81.520000 234.780000 82.070000 234.920000 ;
      RECT 80.760000 234.780000 81.310000 234.920000 ;
      RECT 80.000000 234.780000 80.550000 234.920000 ;
      RECT 79.240000 234.780000 79.790000 234.920000 ;
      RECT 78.480000 234.780000 79.030000 234.920000 ;
      RECT 77.720000 234.780000 78.270000 234.920000 ;
      RECT 76.960000 234.780000 77.510000 234.920000 ;
      RECT 76.200000 234.780000 76.750000 234.920000 ;
      RECT 75.440000 234.780000 75.990000 234.920000 ;
      RECT 74.680000 234.780000 75.230000 234.920000 ;
      RECT 73.920000 234.780000 74.470000 234.920000 ;
      RECT 73.160000 234.780000 73.710000 234.920000 ;
      RECT 72.400000 234.780000 72.950000 234.920000 ;
      RECT 71.640000 234.780000 72.190000 234.920000 ;
      RECT 70.880000 234.780000 71.430000 234.920000 ;
      RECT 70.120000 234.780000 70.670000 234.920000 ;
      RECT 69.360000 234.780000 69.910000 234.920000 ;
      RECT 68.600000 234.780000 69.150000 234.920000 ;
      RECT 67.840000 234.780000 68.390000 234.920000 ;
      RECT 67.080000 234.780000 67.630000 234.920000 ;
      RECT 66.320000 234.780000 66.870000 234.920000 ;
      RECT 65.560000 234.780000 66.110000 234.920000 ;
      RECT 64.800000 234.780000 65.350000 234.920000 ;
      RECT 64.040000 234.780000 64.590000 234.920000 ;
      RECT 63.280000 234.780000 63.830000 234.920000 ;
      RECT 62.520000 234.780000 63.070000 234.920000 ;
      RECT 61.760000 234.780000 62.310000 234.920000 ;
      RECT 61.000000 234.780000 61.550000 234.920000 ;
      RECT 60.240000 234.780000 60.790000 234.920000 ;
      RECT 59.480000 234.780000 60.030000 234.920000 ;
      RECT 58.720000 234.780000 59.270000 234.920000 ;
      RECT 57.960000 234.780000 58.510000 234.920000 ;
      RECT 57.200000 234.780000 57.750000 234.920000 ;
      RECT 56.440000 234.780000 56.990000 234.920000 ;
      RECT 55.680000 234.780000 56.230000 234.920000 ;
      RECT 54.920000 234.780000 55.470000 234.920000 ;
      RECT 54.160000 234.780000 54.710000 234.920000 ;
      RECT 53.400000 234.780000 53.950000 234.920000 ;
      RECT 52.640000 234.780000 53.190000 234.920000 ;
      RECT 51.880000 234.780000 52.430000 234.920000 ;
      RECT 51.120000 234.780000 51.670000 234.920000 ;
      RECT 50.360000 234.780000 50.910000 234.920000 ;
      RECT 49.600000 234.780000 50.150000 234.920000 ;
      RECT 48.840000 234.780000 49.390000 234.920000 ;
      RECT 48.080000 234.780000 48.630000 234.920000 ;
      RECT 47.320000 234.780000 47.870000 234.920000 ;
      RECT 46.560000 234.780000 47.110000 234.920000 ;
      RECT 45.800000 234.780000 46.350000 234.920000 ;
      RECT 45.040000 234.780000 45.590000 234.920000 ;
      RECT 44.280000 234.780000 44.830000 234.920000 ;
      RECT 43.520000 234.780000 44.070000 234.920000 ;
      RECT 42.760000 234.780000 43.310000 234.920000 ;
      RECT 42.000000 234.780000 42.550000 234.920000 ;
      RECT 41.240000 234.780000 41.790000 234.920000 ;
      RECT 40.480000 234.780000 41.030000 234.920000 ;
      RECT 39.720000 234.780000 40.270000 234.920000 ;
      RECT 38.960000 234.780000 39.510000 234.920000 ;
      RECT 38.200000 234.780000 38.750000 234.920000 ;
      RECT 37.440000 234.780000 37.990000 234.920000 ;
      RECT 36.680000 234.780000 37.230000 234.920000 ;
      RECT 35.920000 234.780000 36.470000 234.920000 ;
      RECT 35.160000 234.780000 35.710000 234.920000 ;
      RECT 34.400000 234.780000 34.950000 234.920000 ;
      RECT 33.640000 234.780000 34.190000 234.920000 ;
      RECT 32.880000 234.780000 33.430000 234.920000 ;
      RECT 32.120000 234.780000 32.670000 234.920000 ;
      RECT 31.360000 234.780000 31.910000 234.920000 ;
      RECT 30.600000 234.780000 31.150000 234.920000 ;
      RECT 29.840000 234.780000 30.390000 234.920000 ;
      RECT 29.080000 234.780000 29.630000 234.920000 ;
      RECT 28.320000 234.780000 28.870000 234.920000 ;
      RECT 27.560000 234.780000 28.110000 234.920000 ;
      RECT 26.800000 234.780000 27.350000 234.920000 ;
      RECT 26.040000 234.780000 26.590000 234.920000 ;
      RECT 25.280000 234.780000 25.830000 234.920000 ;
      RECT 24.520000 234.780000 25.070000 234.920000 ;
      RECT 23.760000 234.780000 24.310000 234.920000 ;
      RECT 23.000000 234.780000 23.550000 234.920000 ;
      RECT 22.240000 234.780000 22.790000 234.920000 ;
      RECT 21.480000 234.780000 22.030000 234.920000 ;
      RECT 20.720000 234.780000 21.270000 234.920000 ;
      RECT 19.960000 234.780000 20.510000 234.920000 ;
      RECT 0.000000 234.780000 19.750000 234.920000 ;
      RECT 0.000000 0.140000 236.930000 234.780000 ;
      RECT 228.200000 0.000000 236.930000 0.140000 ;
      RECT 226.490000 0.000000 227.990000 0.140000 ;
      RECT 224.780000 0.000000 226.280000 0.140000 ;
      RECT 223.070000 0.000000 224.570000 0.140000 ;
      RECT 221.360000 0.000000 222.860000 0.140000 ;
      RECT 219.650000 0.000000 221.150000 0.140000 ;
      RECT 217.940000 0.000000 219.440000 0.140000 ;
      RECT 216.230000 0.000000 217.730000 0.140000 ;
      RECT 214.520000 0.000000 216.020000 0.140000 ;
      RECT 212.810000 0.000000 214.310000 0.140000 ;
      RECT 211.100000 0.000000 212.600000 0.140000 ;
      RECT 209.390000 0.000000 210.890000 0.140000 ;
      RECT 207.680000 0.000000 209.180000 0.140000 ;
      RECT 205.970000 0.000000 207.470000 0.140000 ;
      RECT 204.260000 0.000000 205.760000 0.140000 ;
      RECT 202.550000 0.000000 204.050000 0.140000 ;
      RECT 200.840000 0.000000 202.340000 0.140000 ;
      RECT 199.130000 0.000000 200.630000 0.140000 ;
      RECT 197.420000 0.000000 198.920000 0.140000 ;
      RECT 195.710000 0.000000 197.210000 0.140000 ;
      RECT 194.000000 0.000000 195.500000 0.140000 ;
      RECT 192.290000 0.000000 193.790000 0.140000 ;
      RECT 190.580000 0.000000 192.080000 0.140000 ;
      RECT 188.870000 0.000000 190.370000 0.140000 ;
      RECT 187.160000 0.000000 188.660000 0.140000 ;
      RECT 185.450000 0.000000 186.950000 0.140000 ;
      RECT 183.740000 0.000000 185.240000 0.140000 ;
      RECT 182.030000 0.000000 183.530000 0.140000 ;
      RECT 180.320000 0.000000 181.820000 0.140000 ;
      RECT 178.610000 0.000000 180.110000 0.140000 ;
      RECT 176.900000 0.000000 178.400000 0.140000 ;
      RECT 175.190000 0.000000 176.690000 0.140000 ;
      RECT 173.480000 0.000000 174.980000 0.140000 ;
      RECT 171.770000 0.000000 173.270000 0.140000 ;
      RECT 170.060000 0.000000 171.560000 0.140000 ;
      RECT 168.350000 0.000000 169.850000 0.140000 ;
      RECT 166.640000 0.000000 168.140000 0.140000 ;
      RECT 164.930000 0.000000 166.430000 0.140000 ;
      RECT 163.220000 0.000000 164.720000 0.140000 ;
      RECT 161.510000 0.000000 163.010000 0.140000 ;
      RECT 159.800000 0.000000 161.300000 0.140000 ;
      RECT 158.090000 0.000000 159.590000 0.140000 ;
      RECT 156.380000 0.000000 157.880000 0.140000 ;
      RECT 154.670000 0.000000 156.170000 0.140000 ;
      RECT 152.960000 0.000000 154.460000 0.140000 ;
      RECT 151.250000 0.000000 152.750000 0.140000 ;
      RECT 149.540000 0.000000 151.040000 0.140000 ;
      RECT 147.830000 0.000000 149.330000 0.140000 ;
      RECT 146.120000 0.000000 147.620000 0.140000 ;
      RECT 144.410000 0.000000 145.910000 0.140000 ;
      RECT 142.700000 0.000000 144.200000 0.140000 ;
      RECT 140.990000 0.000000 142.490000 0.140000 ;
      RECT 139.280000 0.000000 140.780000 0.140000 ;
      RECT 137.570000 0.000000 139.070000 0.140000 ;
      RECT 135.860000 0.000000 137.360000 0.140000 ;
      RECT 134.150000 0.000000 135.650000 0.140000 ;
      RECT 132.440000 0.000000 133.940000 0.140000 ;
      RECT 130.730000 0.000000 132.230000 0.140000 ;
      RECT 129.020000 0.000000 130.520000 0.140000 ;
      RECT 127.310000 0.000000 128.810000 0.140000 ;
      RECT 125.600000 0.000000 127.100000 0.140000 ;
      RECT 123.890000 0.000000 125.390000 0.140000 ;
      RECT 122.180000 0.000000 123.680000 0.140000 ;
      RECT 120.470000 0.000000 121.970000 0.140000 ;
      RECT 118.760000 0.000000 120.260000 0.140000 ;
      RECT 117.050000 0.000000 118.550000 0.140000 ;
      RECT 115.340000 0.000000 116.840000 0.140000 ;
      RECT 113.630000 0.000000 115.130000 0.140000 ;
      RECT 111.920000 0.000000 113.420000 0.140000 ;
      RECT 110.210000 0.000000 111.710000 0.140000 ;
      RECT 108.500000 0.000000 110.000000 0.140000 ;
      RECT 106.790000 0.000000 108.290000 0.140000 ;
      RECT 105.080000 0.000000 106.580000 0.140000 ;
      RECT 103.370000 0.000000 104.870000 0.140000 ;
      RECT 101.660000 0.000000 103.160000 0.140000 ;
      RECT 99.950000 0.000000 101.450000 0.140000 ;
      RECT 98.240000 0.000000 99.740000 0.140000 ;
      RECT 96.530000 0.000000 98.030000 0.140000 ;
      RECT 94.820000 0.000000 96.320000 0.140000 ;
      RECT 93.110000 0.000000 94.610000 0.140000 ;
      RECT 91.400000 0.000000 92.900000 0.140000 ;
      RECT 89.690000 0.000000 91.190000 0.140000 ;
      RECT 87.980000 0.000000 89.480000 0.140000 ;
      RECT 86.270000 0.000000 87.770000 0.140000 ;
      RECT 84.560000 0.000000 86.060000 0.140000 ;
      RECT 82.850000 0.000000 84.350000 0.140000 ;
      RECT 81.140000 0.000000 82.640000 0.140000 ;
      RECT 79.430000 0.000000 80.930000 0.140000 ;
      RECT 77.720000 0.000000 79.220000 0.140000 ;
      RECT 76.010000 0.000000 77.510000 0.140000 ;
      RECT 74.300000 0.000000 75.800000 0.140000 ;
      RECT 72.590000 0.000000 74.090000 0.140000 ;
      RECT 70.880000 0.000000 72.380000 0.140000 ;
      RECT 69.170000 0.000000 70.670000 0.140000 ;
      RECT 67.460000 0.000000 68.960000 0.140000 ;
      RECT 65.750000 0.000000 67.250000 0.140000 ;
      RECT 64.040000 0.000000 65.540000 0.140000 ;
      RECT 62.330000 0.000000 63.830000 0.140000 ;
      RECT 60.620000 0.000000 62.120000 0.140000 ;
      RECT 58.910000 0.000000 60.410000 0.140000 ;
      RECT 57.200000 0.000000 58.700000 0.140000 ;
      RECT 55.490000 0.000000 56.990000 0.140000 ;
      RECT 53.780000 0.000000 55.280000 0.140000 ;
      RECT 52.070000 0.000000 53.570000 0.140000 ;
      RECT 50.360000 0.000000 51.860000 0.140000 ;
      RECT 48.650000 0.000000 50.150000 0.140000 ;
      RECT 46.940000 0.000000 48.440000 0.140000 ;
      RECT 45.230000 0.000000 46.730000 0.140000 ;
      RECT 43.520000 0.000000 45.020000 0.140000 ;
      RECT 41.810000 0.000000 43.310000 0.140000 ;
      RECT 40.100000 0.000000 41.600000 0.140000 ;
      RECT 38.390000 0.000000 39.890000 0.140000 ;
      RECT 36.680000 0.000000 38.180000 0.140000 ;
      RECT 34.970000 0.000000 36.470000 0.140000 ;
      RECT 33.260000 0.000000 34.760000 0.140000 ;
      RECT 31.550000 0.000000 33.050000 0.140000 ;
      RECT 29.840000 0.000000 31.340000 0.140000 ;
      RECT 28.130000 0.000000 29.630000 0.140000 ;
      RECT 26.420000 0.000000 27.920000 0.140000 ;
      RECT 24.710000 0.000000 26.210000 0.140000 ;
      RECT 23.000000 0.000000 24.500000 0.140000 ;
      RECT 21.290000 0.000000 22.790000 0.140000 ;
      RECT 19.580000 0.000000 21.080000 0.140000 ;
      RECT 17.870000 0.000000 19.370000 0.140000 ;
      RECT 16.160000 0.000000 17.660000 0.140000 ;
      RECT 14.450000 0.000000 15.950000 0.140000 ;
      RECT 12.740000 0.000000 14.240000 0.140000 ;
      RECT 11.030000 0.000000 12.530000 0.140000 ;
      RECT 9.320000 0.000000 10.820000 0.140000 ;
      RECT 0.000000 0.000000 9.110000 0.140000 ;
    LAYER metal3 ;
      RECT 0.000000 0.000000 236.930000 234.920000 ;
    LAYER metal4 ;
      RECT 0.000000 0.000000 236.930000 234.920000 ;
    LAYER metal5 ;
      RECT 0.000000 0.000000 236.930000 234.920000 ;
    LAYER metal6 ;
      RECT 0.000000 0.000000 236.930000 234.920000 ;
    LAYER metal7 ;
      RECT 0.000000 0.000000 236.930000 234.920000 ;
    LAYER metal8 ;
      RECT 0.000000 0.000000 236.930000 234.920000 ;
    LAYER metal9 ;
      RECT 0.000000 0.000000 236.930000 234.920000 ;
    LAYER metal10 ;
      RECT 0.000000 0.000000 236.930000 234.920000 ;
  END
END aes128key

END LIBRARY
